��  CCircuit��  CPart          ���  CRailEnd�� 	 CTerminal  �0�1           �          �,�4 	    ��  �P�Q           �          �L�T     �� 
 CResistorH��  CValue  H�h�10k        ��@      �?k �  8�M�           �        �  d�y�           �          L�d�     ��  Hnh|10k        ��@      �?k �  8�M�           �        �  d�y�           �          L|d�     ��  H>hL10k        ��@      �?k �  8PMQ                     �  dPyQ           �          LLdT     �� 	 CPushMake��  CKey  � ��   �  � �� �           �        �  ��           �          � ��     ��  � Xt    �  � P� Q           �        �  PQ                      � HT "    ��  � ��  $ �  � �� �           �        �  ��           �          � x� &              ���  CWire  � 0� Q )�  � 0�1 )�  xP�Q )�  x�y� )�  xPy� )�  �9� )�  �9� )�  P9Q  )�  � �� � )�  � P� �           �                      + 	   ,    /     -   0     .   1     .   2     /   3 "   # 1   3 &   ' 0 + " * 	     , -   '  #  &  * 2             � ��         @         