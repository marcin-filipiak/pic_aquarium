��  CCircuit��  CPart          ���  CPot��  CValue  � �� �45k          ��@      �?k ��  CSlider  � ��  �� 	 CTerminal  � �� �     �*�q@͝_\�f)?�  � �� �    �������=        �  ��    �������=͝_\�f)�  � ��   
 ��  CEarth�  ��     �������=Ν_\�f)?  �$     ��  CRailEnd�  0�E�    �*�q@          D�L�     ��  CVPos�  � 9� G5V'          @      �? V�  � @� A    ������@   ��f)�  � <� D     �� 	 CResistor�  � a� o3.3k          ȩ@      �?k �  � H� ]     ������@ʝ_\�f)?�  � t� �    �*�q@ʝ_\�f)�  � \� t               ���  CWire  ��  �  � �1�  �  � �� �  �  � @� I  �  � @� A           �                      "          !   !    "     %   $     #   #    %   $            � ��         @         